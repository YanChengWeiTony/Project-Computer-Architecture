module Instruction_Memory
(
    addr_i, 
    data_o
);

// Ports
input   [31:0]		addr_i;
output  [31:0]      data_o;

// Instruction memory
reg     [31:0]		memory 	[0:255];

assign  data_o = memory[addr_i>>2];  

endmodule